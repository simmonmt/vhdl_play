package libbase is
  function log2ceil(x: natural) return integer;
end libbase;
